library verilog;
use verilog.vl_types.all;
entity SineWaveGenerator_vlg_vec_tst is
end SineWaveGenerator_vlg_vec_tst;
