library verilog;
use verilog.vl_types.all;
entity SineWave_vlg_vec_tst is
end SineWave_vlg_vec_tst;
