library verilog;
use verilog.vl_types.all;
entity driverSPWMGenerator_vlg_vec_tst is
end driverSPWMGenerator_vlg_vec_tst;
